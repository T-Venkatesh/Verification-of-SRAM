`ifndef _bp_
`define _bp_

class basepkt;
rand bit[7:0]data_in;
randc bit[5:0]addr;
bit en;
bit wr;
bit [7:0]data_out;
endclass
`endif   
